ecc_curve_iram/ecc_vars.vhd