ecc_fp_dram/ecc_fp_dram_sh.vhd